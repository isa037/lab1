
library ieee;
use ieee.numeric_std.all;



package pkg is
  type array8 is array (natural range <>) of signed(7 downto 0);
end package;

package body pkg is
	

end package body;
