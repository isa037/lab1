LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--use ieee.fixed_pkg.all;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MULTIPLIER IS
	GENERIC ( N, M : INTEGER:=24);
	PORT (	A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			B : IN signed(M-1 DOWNTO 0);
			OUTPUT :	OUT STD_LOGIC_VECTOR(M+N-1 DOWNTO 0));
END MULTIPLIER;

ARCHITECTURE BEHAVIOR OF MULTIPLIER IS
BEGIN	

	OUTPUT<=std_logic_vector(to_signed(A)*B);

END BEHAVIOR;
