LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--use ieee.fixed_pkg.all;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MULTIPLIER IS
	GENERIC ( N, M, K : INTEGER:=24);
	PORT (	A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			B : IN signed(M-1 DOWNTO 0);
			OUTPUT :	OUT STD_LOGIC_VECTOR(K-1 DOWNTO 0));
END MULTIPLIER;

ARCHITECTURE BEHAVIOR OF MULTIPLIER IS
	
	signal OUTPUT_tmp : std_logic_vector(N+M-1 downto 0);
	
BEGIN	

	OUTPUT_tmp<=std_logic_vector(signed(A)*B);
	OUTPUT<=OUTPUT_tmp(N+M-1 downto N+M-K);

END BEHAVIOR;
