LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--use ieee.fixed_pkg.all;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ADDER IS
	GENERIC ( N : INTEGER:=9);
	PORT (	A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			B : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			OUTPUT :	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END ADDER;

ARCHITECTURE BEHAVIOR OF ADDER IS
BEGIN	

	OUTPUT<=std_logic_vector(signed(A)+signed(B));

END BEHAVIOR;
